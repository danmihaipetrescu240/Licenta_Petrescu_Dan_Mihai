module dense_layer1(
    input clock,
    input enable,
    input reset,
    input signed [15:0] imagine_trasa [0:195],
    output signed [15:0] iesire_layer [0:31],
    output layer_terminat
    );
    
    reg signed [31:0] dense1_retea [0:31];
    reg signed [15:0] relu_retea [0:31];
localparam signed [7:0] VECTOR_BIASURI_LAYER2 [0:31] = '{ 12, 4, -6, 20, 6, 13, -4, 7, 6, 8, 8, 19, 18, 10, -7, 18, 6, -13, 4, 10, -2, -11, 14, 1, -6, 3, -18, 12, 23, 10, -8, -1 };
  
  localparam signed [7:0] VECTOR_WEIGHTS_LAYER2 [0:31] [0:195] = '{
{ 3, -1, 7, 24, 19, 29, 12, 1, 22, 31, 15, 6, -3, 7, -8, 9, 21, 52, 56, 44, 24, -2, -14, 10, 19, 4, 20, 18, 7, 36, 33, 9, 12, 8, 17, -2, 1, 3, -11, -8, -10, -11, 18, 23, 24, 1, -6, 7, 9, 2, -11, -10, -2, -2, 24, 31, 27, 15, 2, -5, -17, -26, -8, 6, -20, -15, -4, 2, 9, 10, 11, 3, -16, -36, -35, -14, 30, 1, -19, -8, -15, -35, 7, 43, -2, 11, 2, 5, 20, 37, 20, -21, -18, -19, -28, -41, -44, 14, 16, 30, 9, 9, 25, 2, -14, -17, -20, -9, -1, 6, 26, 22, 12, 42, -9, -46, -43, -25, -27, -6, 3, 11, 14, 22, 22, 28, 23, 33, -18, -21, -30, -29, -9, 13, 24, 13, 8, 14, -4, 1, 5, 24, -7, 10, 21, 14, 26, 28, 9, 12, 0, 22, 13, 32, 1, 49, 27, 7, 29, 32, 15, 9, -7, 3, -9, 13, -15, 22, 7, 26, 12, 17, 16, 14, 9, 13, 3, -6, -4, 4, 20, 18, -3, -1, -26, -19, -20, 9, 1, -29, -25, 0, 7, 18, -1, 5 },
{ 1, 6, 13, 11, 26, 46, 43, 21, 22, 34, 12, 16, -8, 6, -8, 6, -10, -4, 12, -7, -4, 3, 10, -1, -10, 10, 0, -4, 4, -37, -34, -16, 18, -4, -8, -5, 2, 1, 4, -14, 5, 20, 12, -32, -21, 2, 13, 4, 7, -19, -14, -15, -4, 14, 2, 4, 23, 13, 4, 15, 10, -3, 10, -8, -5, 2, -2, 16, 9, 29, 31, -25, 0, 23, 23, 14, 8, -11, -7, 5, 3, 13, 5, 2, 7, 15, 5, 15, 14, -15, -11, -10, -14, -8, 7, 9, 55, -4, 14, 26, 2, -23, -59, -29, 11, 8, -7, -15, -22, -9, 24, 26, 8, 12, -43, -73, -63, 27, 41, 12, -4, -8, -17, -12, 26, 4, -2, -31, -82, -50, -1, 47, 43, -2, -1, 2, -11, -8, 17, 15, 14, -21, -40, -1, -2, 24, 29, 5, 3, 10, -5, -7, -5, 4, 2, -11, 0, -10, -6, 3, 21, 15, -5, 0, 1, -7, -7, -22, 5, -29, -20, -12, -9, 0, 9, 6, 2, 1, -12, -18, 9, 5, -9, -12, -20, -6, 2, -6, -25, -23, -37, -23, -16, 17, 5, -8 },
{ 5, -4, -7, -4, -24, -47, -37, -1, 19, -31, -22, 1, -9, 3, 3, 0, 12, 5, 32, 33, 34, 20, 16, 4, -2, -23, 8, -1, 11, 25, 24, 24, 16, 26, 20, 28, 28, 26, 5, -17, -11, 3, 23, 1, -1, -16, 1, -1, 21, 20, 16, 11, 4, -18, -52, -14, -13, 15, -2, -5, -7, -14, -20, -14, 11, 18, 5, -9, -127, -12, -24, 24, -7, -16, -32, -25, -36, -12, 5, 28, 18, 3, -71, -6, -37, 16, -24, -26, -2, -2, 8, 10, -7, 10, 21, -25, -30, 21, 6, 13, 4, 11, -11, -22, 6, 4, 0, 5, 4, -12, -1, 27, 28, 41, 33, -2, -30, -26, -15, -12, 2, 7, 3, 0, 6, 11, -20, 29, 24, 8, -12, 3, -4, 4, 17, 8, 3, -14, -8, 20, -12, 38, 14, 15, 11, 1, -2, 1, 20, 13, 3, -20, 1, 15, 7, 48, -8, 7, 2, 18, 9, 6, 6, 13, 7, 19, 22, 6, 5, 6, 6, 16, 7, 13, 16, 13, 17, 11, 24, 34, 43, 6, -7, 13, 23, -7, -4, 9, 18, 17, 18, 17, 31, 17, 8, 8 },
{ 4, -5, 2, -3, -13, -8, -10, 10, -13, -22, -3, 0, 6, -4, -8, 13, 2, 6, -27, -31, 5, 3, -2, 0, 8, 3, -29, -7, 0, 14, 22, 5, -23, -2, 8, 11, 7, -9, -14, -1, 16, -6, 5, -14, -7, -20, -10, 4, 4, -1, -5, -4, -2, 0, 10, 32, -36, -12, -27, -21, 0, 7, 10, -3, -3, 6, 13, 1, 34, 35, 1, -35, -38, -27, 4, 0, 9, -3, -17, -2, 0, 32, 61, 46, -13, -34, -19, -23, 0, 19, 39, 10, 1, -6, -12, -26, -13, 2, 6, -16, -32, -58, -4, 24, 41, 26, 5, -2, -15, -30, -36, -35, 20, -1, -19, -61, -81, -27, 12, 20, 8, -7, -9, -39, -45, -19, -20, 15, 17, -14, -48, -52, -30, 3, 9, -4, -6, -41, -19, 13, 13, -6, 22, 24, 10, -3, -16, 5, 10, -2, -20, -13, -11, 8, 7, 17, 26, 11, 7, 14, 1, -1, -9, -19, -34, -39, -15, 27, 6, 36, 19, 1, 23, 24, 6, 2, -6, -36, -10, 13, 8, -4, 8, 5, 17, -2, -21, 9, -15, -3, 10, 18, 26, 18, -7, 7 },
{ -7, -8, -7, 0, 7, 4, 2, 27, 33, 0, -8, -1, 6, 0, -8, 13, 6, -24, 15, 17, 33, 26, 19, -12, -13, -4, 5, 3, 0, 9, -33, -10, -2, 9, 15, 21, 28, 19, 4, -16, -12, 11, 4, -16, -23, -28, -27, 6, -2, 6, 27, 40, 30, 22, -25, -18, 13, 5, -12, -28, -15, -11, 2, 7, 39, 33, 25, 38, 34, 7, 8, -8, -35, -3, -9, -10, -6, 1, -14, -1, 17, 27, 29, 5, 1, -15, -15, 4, 5, 8, 12, -24, -42, -12, -3, 11, 9, 1, -22, -7, 25, 16, 3, 13, 16, -19, -33, -24, -4, 10, 7, 28, -19, -3, 25, 17, 8, 8, -32, -21, 2, -32, -20, 1, 21, 26, 24, -23, 0, 11, 17, -8, -27, -5, -5, -27, -13, 14, 19, 20, 23, 17, 33, 20, 10, 2, 7, -3, 8, -15, 0, 21, -17, -1, -2, 43, 9, 22, 22, 22, 17, 5, 7, 8, -6, 27, 6, -23, 3, 2, -8, -3, 27, 31, 32, 16, 22, 21, 21, 16, 20, -4, -5, -3, -17, -16, 15, 28, 11, -9, -8, -1, -17, 15, -8, 9 },
{ 9, 6, 4, -11, -25, -24, -27, 3, -63, -34, -37, -2, -6, 2, -7, 1, -5, -24, -36, -36, -22, -5, 7, -4, 7, -16, -3, -12, 5, 9, -13, -1, -17, 4, -5, -6, -11, -12, -8, -2, 18, 7, 14, 26, 0, 7, 1, 3, 15, 8, 15, 8, 4, 13, 21, 22, 9, -6, -10, 16, 2, 7, 20, 30, 23, 22, 23, 24, 58, 36, 17, 8, 5, 19, 6, 26, 37, 35, 16, 18, 8, 8, 50, 72, 18, 22, 6, 13, 0, -2, 11, 12, 5, 8, -7, -36, -29, 29, 5, -14, 0, -3, -9, -7, -30, -14, -5, 2, -2, -5, -6, -44, 2, -17, -3, 0, 0, -15, -29, -8, -1, 3, 2, -1, -3, -27, 25, 0, 5, 10, 9, 2, 3, 1, -1, 4, 5, 4, 4, -30, -5, -27, -9, 6, 3, -8, -4, -14, -1, -11, -10, -4, 3, -29, 5, -30, -7, -4, -1, 3, -8, 2, 1, -19, -9, -10, -6, -25, -6, 34, 26, 17, 13, 20, 16, 13, 16, 12, 5, 8, 4, -18, 7, 0, -17, 1, 46, 53, 60, 63, 70, 69, 48, 27, -6, 7 },
{ 7, -2, 3, 3, 12, 33, 8, -2, -28, 20, 25, 29, -5, 7, 1, -7, -23, -1, -10, 0, -57, -56, -41, -10, 16, 8, 9, -1, 11, 20, 6, 3, -5, -18, -51, -21, 3, 14, 3, 0, -18, -20, 24, 19, 5, 5, 4, -10, -37, -11, 17, 20, 14, -3, -9, -3, 37, 17, -1, 4, 3, 1, -51, 1, 34, 18, -7, -21, -40, -5, 39, 37, 9, -11, 1, -48, -56, 34, 30, -3, -4, -10, -21, 4, 26, 9, 1, -16, -36, -17, 24, 22, 10, 8, 0, -16, -40, -18, 14, -14, 7, -34, -3, 20, 24, 8, 10, 4, 21, -41, -52, -22, 34, -14, 2, -5, 5, 20, 36, 5, 3, 33, 0, -50, -60, 5, 23, 15, 4, -17, -12, -2, 13, -5, 10, 1, -23, -52, -66, 10, 13, 3, 6, 4, 4, -9, 2, 5, -7, -24, -10, -35, -39, 17, 4, -11, 26, 21, 3, 3, 0, 4, -8, -22, -10, -7, -28, 27, 7, 22, 17, 5, -15, -7, 6, -18, -15, -7, -26, -21, -25, 4, -9, -14, -29, -28, -40, -9, -46, -55, -29, -41, -42, -28, 6, -2 },
{ -6, 2, 1, 28, 28, 45, 19, 2, 58, 28, 36, 23, -6, -3, -3, 28, 22, 45, 65, 65, 39, 25, 16, 38, 24, 51, 41, 13, -8, 12, 9, 4, 0, 15, 4, 9, 16, 16, 10, -15, 9, 44, -9, -18, -2, -10, 1, 14, 6, 6, 7, -6, -15, -19, 14, 6, -40, -10, 8, 8, 11, -2, -1, -1, -8, -14, -8, -11, -12, 3, -35, -1, 27, 18, -5, -14, -3, 11, -14, 2, 9, 22, 40, 14, -32, -4, 26, 0, -18, -27, 28, 24, 1, -4, 1, 15, 30, 18, -25, 7, 5, 3, -21, 8, 37, 14, 7, 10, 9, -16, 11, 33, -11, 9, 17, 0, -4, 14, 20, -3, 3, 11, -5, -2, 11, 22, -23, -16, -3, 25, 7, 11, 2, 5, 24, 23, -5, 16, 24, 6, -15, 13, 13, 21, 22, 19, 16, 22, 15, 15, 3, 19, 11, -14, 3, 47, 1, -17, 2, 8, 24, 0, 4, -1, 6, 13, 11, -30, 5, -7, -15, -7, -8, -2, 0, -3, 14, 19, 20, 8, 25, 1, -2, 18, 25, 1, 7, 19, 25, 15, 4, 10, 32, -3, 12, 3 },
{ 3, 3, -6, 12, 2, 0, 4, 15, 42, 11, 8, 4, 7, 5, 2, 2, 7, 17, 45, 31, 27, 9, -7, 16, 2, -13, 8, 10, -9, -2, -19, 4, 14, 16, 10, 14, 8, -1, 1, 15, -10, 4, 16, -5, -26, -1, 8, 18, 26, 40, 33, 25, 15, 18, 9, 6, 12, -11, -13, -19, 2, 10, 15, 36, 38, 25, 0, 10, -7, 6, 25, 2, -25, -7, -11, -22, -42, -49, -35, -23, -22, -19, -15, 34, 14, -6, -27, -25, -15, -21, -28, -34, -35, -13, -23, -37, -37, 16, -1, -3, -27, 5, -6, -2, 10, -1, -15, -28, -18, -40, -13, 29, -18, 2, -2, -16, 2, 6, 11, -7, -17, -33, -15, -22, 2, 42, 9, -7, -5, -16, -13, -17, -7, -15, 4, 4, 9, -5, 23, 41, 12, 40, 5, -5, 6, 8, 31, 25, 26, 30, 35, 23, 28, 48, -7, 38, 18, 4, 1, 27, 21, 29, 28, 31, 20, 35, 22, 4, 6, 0, -11, 4, 26, 26, 36, 34, 20, 33, 13, 8, 35, 15, 8, -5, -15, -17, 3, 13, 16, 21, 39, 21, -11, -24, 16, -1 },
{ -3, -3, 10, -9, 10, 4, 9, 19, -31, 14, 1, -17, -8, -2, -7, 1, -15, -43, -29, -46, -17, -12, 1, -5, -20, 17, -9, -7, -4, -16, -13, 13, -11, -19, -3, -5, -8, -13, -10, -13, 3, 3, -21, 2, -6, -10, 6, 6, 5, 14, 10, 3, 9, -9, -3, -8, -5, 4, -9, 16, 18, -2, 3, 14, -7, 8, -8, -8, -7, 7, 13, -15, 0, 9, 3, 13, 22, 29, -17, 2, 3, 6, -21, -6, 19, 24, 22, 13, 4, 2, -1, 20, 12, 4, 17, 29, -17, -25, -6, 12, 0, -18, -12, 10, 2, 11, 3, 7, -11, -29, -45, -54, -2, -22, -33, -25, 14, -1, 0, 22, 16, -7, -12, -27, -26, -12, 16, -60, -74, -24, 9, -1, 5, 8, -1, -5, -6, -38, -17, 13, -5, -57, -26, -14, -10, -17, -2, -1, -9, -13, -13, -32, -4, -8, -5, -49, 0, 4, -1, -3, 5, 4, 8, -2, -16, -11, -7, -32, 1, -20, -8, -4, -1, 1, -6, 4, -2, 8, 6, -11, -13, -9, -1, 9, 5, 24, 37, 16, 12, 38, 14, 25, 23, 20, 3, -9 },
{ 9, 9, 1, -6, 27, 0, 12, -7, -26, -10, -24, -24, 7, -8, -7, -2, 8, -1, -9, 8, -5, 14, 6, 7, 20, 28, -4, 14, -6, 2, -28, -25, -2, 12, -5, -13, -5, -4, 11, 15, 53, 20, -6, -33, -31, -33, -1, -9, -16, 7, -2, -7, 6, 14, 49, 73, -14, -22, -23, 2, 10, -16, -15, -9, -2, 2, 15, 8, 66, 26, -31, -31, -6, 18, 32, 5, -45, -41, -27, -18, -18, -3, 44, 22, -21, -20, -7, 18, 30, 32, 2, -13, -12, 6, -7, -16, -23, -39, -1, -3, 3, 15, 19, 24, 13, 6, 20, 4, -21, -24, -30, -14, -7, -3, 2, 8, 15, 14, 34, 1, 16, -9, -13, -18, -7, -25, -8, -6, -3, 25, 7, 16, 19, 4, -5, -3, -9, -13, -1, -20, -14, 8, -41, -29, -14, -12, 1, 1, 8, 3, 9, 25, 14, -7, -3, 12, -34, -59, -23, -5, 7, 7, 5, 10, 26, 46, 24, -3, -7, 5, -8, -12, -14, -1, -3, 11, 23, 24, 32, 47, 21, -12, 7, 11, 21, 15, 4, 12, 13, 2, -7, -23, -1, -5, -12, 7 },
{ 9, -6, 3, 11, 23, 30, 30, -16, 11, 34, 29, 22, -1, 6, 5, -1, 13, 5, 30, 11, -18, -6, -8, 5, 18, 13, 17, 19, -3, -5, -2, -24, -22, -25, -24, -16, -11, -1, -3, 3, 1, 1, -11, 15, 8, -12, -8, -36, -19, -5, -8, -9, -8, -2, 11, 19, 2, -11, -20, -6, -19, -23, -4, 0, -6, -10, -3, -18, 14, -21, 9, -10, -30, -7, -12, 2, 12, -3, -1, -11, -20, 1, 23, 1, 0, -42, -34, 3, 2, 32, 35, -6, -2, -3, -15, -13, 2, -12, 17, 9, 4, 21, 15, 41, 13, -3, 24, 18, -14, 16, 38, 1, -21, 12, 6, 15, 15, 20, -9, 15, 46, 30, 16, 17, 10, -9, -19, 10, 12, 15, 9, 7, 2, 28, 28, 15, 6, -8, 7, -18, 17, 24, -4, -4, 4, 5, 8, -8, -11, -14, 3, -5, -18, 4, 2, 16, 2, -15, -8, -7, -14, -32, -17, -28, -20, -21, -7, 16, -1, 3, -7, -22, -26, -32, -36, -24, -23, -6, -11, 5, 17, -1, 5, -19, -13, -38, -69, -61, -40, -55, -29, -27, -31, -12, -16, -8 },
{ 4, -5, -1, -3, -8, -21, -14, -13, -31, -20, -33, -8, 0, 0, -3, -5, -8, -18, -28, -38, -61, -67, -61, -27, -23, -24, -26, -3, 0, -11, -5, -10, -14, -41, -18, -26, -24, -19, 2, -3, 4, -23, -26, 8, 1, -14, -29, -7, 4, 5, 16, 18, 28, 17, -4, 23, -18, -16, 5, -7, -19, -17, 19, 16, -4, 1, 6, -2, 10, 2, -5, -16, -22, -25, -16, 3, 32, 25, 5, -28, -19, -10, 11, 11, 11, 5, -9, -2, 0, 13, -9, 24, 21, -24, -9, -15, 14, 12, 1, 5, 1, -17, -8, -2, -9, 28, 27, -12, -8, 6, -8, -31, 8, -15, -10, 8, 1, 5, 7, 19, -11, -34, -1, 6, -7, 8, 20, -26, -25, -12, -9, 8, 17, -18, -44, -28, -23, -29, 2, 31, -7, -28, -23, -16, 3, 2, 2, -14, -5, -29, -23, -26, 26, -6, -3, -33, 1, -3, 13, 11, 14, 11, 8, -11, 1, 9, -6, 5, -5, -23, -18, -14, -17, -12, -13, 1, -13, 6, 2, 15, 15, 7, 1, 10, 5, 14, 32, -6, 1, 18, 4, 11, 11, 21, 8, 5 },
{ 6, -6, -9, -20, -25, -36, -28, -31, -19, -28, -28, -19, 1, -7, 0, -4, -7, -55, -74, -76, -112, -79, -29, 7, 8, 5, 8, -7, 10, 13, -10, -4, -18, -18, -15, -30, -10, 0, -4, 10, 23, 5, 19, 18, 7, 8, 15, 17, 13, 14, 18, 12, 10, 7, 9, 18, -5, 16, 18, 18, 26, 11, -2, 3, 3, 9, 16, 13, 21, 11, -23, 19, 12, 19, 23, 3, -26, -35, -9, -9, 1, 2, 6, 23, 7, 7, 24, 15, 20, 24, 3, 2, 0, -3, 21, 13, -2, 9, 12, 29, 3, 15, 31, 27, 30, 17, 19, 12, 5, 2, -30, -15, 13, -12, -25, -18, 3, 13, 35, 17, 23, -3, 1, 7, -30, -22, -18, 10, -26, -38, -64, -39, -28, -9, -9, -15, -2, -18, -36, 0, 8, 0, -14, -37, -30, -41, -14, -14, -12, -16, 8, -2, -5, -13, -10, 20, 6, 10, 7, 5, 1, -2, -19, 6, -5, 9, -8, 5, 7, 28, 30, 32, 22, 49, 30, 15, 19, 7, 9, 20, -33, -24, 4, -2, 31, 42, 47, 56, 51, 40, 44, 17, 8, 17, -1, 6 },
{ 2, -6, 10, -4, 9, 6, 27, 24, -9, 21, 6, -1, -8, -3, 5, 6, -13, -9, -18, 2, -9, 1, 11, 0, -18, 10, -5, -14, -1, 0, -7, -6, -4, -6, -2, 5, 11, 21, 19, 8, -14, -41, -9, -3, 5, 0, -20, 12, 14, 1, 7, 24, 20, 6, -28, -67, 13, 3, 8, 12, 0, -2, 2, -9, 6, 32, 28, 2, -15, -61, 15, 15, 5, 0, 6, -11, -17, -50, 3, 11, 20, 10, -15, -73, -15, 8, 14, 21, 1, -16, -46, -52, -22, -14, 1, 19, 15, -41, 10, -6, 19, 22, 16, -26, -30, -26, -29, -5, 21, 17, 13, -12, 2, -8, 9, 30, 30, 0, -5, -14, -9, 21, 23, 16, -11, -10, 14, 5, -6, 12, 33, 31, -12, -14, 22, 22, 18, -3, -6, -13, 13, 18, 14, 14, 11, 19, 4, 1, 24, 10, 4, -1, 8, 2, -10, -19, 5, 19, 7, 6, 10, 20, 13, 4, 8, 10, -2, -18, -4, 12, 9, 2, -6, 6, -5, -9, -16, -27, 0, 13, -13, 8, -8, -4, 25, 26, -3, -35, -17, -30, -73, -30, 6, -7, 5, 3 },
{ -3, -2, -7, -10, -12, 0, -10, -3, -6, -34, -35, -1, 8, -3, 4, 10, -4, -34, -16, -36, -37, -30, -21, -34, -17, -23, -3, 24, 0, -13, -29, -34, -33, -26, -30, -46, -49, -36, -34, -31, -8, -3, 1, 30, -27, -14, -4, -2, 13, 11, 15, 8, 3, -7, -4, 11, 35, -1, -18, -21, -4, 20, 28, 31, 28, 35, 12, 22, 42, 18, 21, 12, 0, 14, 16, 19, 28, 16, 14, 11, 19, 13, 57, 67, 20, 30, 14, 5, -2, 11, 10, -7, -20, -14, -21, -24, -34, 56, 8, 0, 7, 6, -1, 1, -7, -27, -10, 7, 5, -4, 26, 21, -19, -13, 14, 1, -12, 7, -6, -11, 23, 10, 1, -3, 12, 23, 29, -30, 3, 5, 2, 0, -1, -3, -4, 6, 4, 18, 6, 4, 20, -27, 2, -19, -17, -23, -5, -20, -9, 0, -7, -1, 10, -4, -5, 10, 0, 4, -8, -3, -11, -21, -18, -29, -29, -1, 25, 5, -6, 28, 33, -1, -3, 1, 2, 12, 13, 12, 14, 16, 19, -12, 1, 4, -5, 5, 22, 47, 59, 71, 66, 59, 66, 41, 10, 3 },
{ 9, -3, 7, 1, 2, 2, -2, 15, 18, 37, 34, 15, 6, -9, -2, 8, 20, 21, -1, -9, 10, 6, 35, 21, 25, 20, 4, -1, 3, 29, 7, 8, -10, 3, -4, 19, 18, 37, 41, 31, 28, 31, 3, -4, 2, 2, -8, -11, 3, 14, 0, 11, 5, 34, 46, 0, -28, 4, -13, -1, 12, 1, 11, 7, 6, -2, -2, 10, 14, 14, -17, -6, -18, -7, -3, -4, 28, 20, -3, 1, -15, 12, 35, 16, -35, -17, -29, -4, -14, -3, 45, 13, -4, -1, -21, -22, 7, -7, 5, -8, -28, -11, -11, -13, 22, 7, -20, -25, -12, -32, 1, -39, 21, 6, 1, -11, -9, 3, 2, -26, -18, -10, -9, 11, -10, -56, -24, 20, 14, 13, -5, -8, -23, -24, 1, 12, 11, 12, -18, -39, 6, -2, 10, 23, 19, 10, 16, 13, 24, 39, 28, 11, -17, -18, 4, 20, 7, 2, 8, 25, 25, 27, 23, 19, 6, -7, -34, 20, 7, 24, 2, 9, 18, 14, 28, 11, 10, -12, -19, -22, -37, -13, 7, 3, 7, -38, -27, -14, -21, -23, -4, -11, -16, -12, -8, 1 },
{ -5, -3, -5, -19, -23, -26, -25, -10, 10, -11, -17, 4, -9, -7, -4, 0, 9, -14, 22, 11, 2, -27, -31, 0, 14, 19, 17, 18, 3, 22, -29, -5, 3, 23, 18, 17, 31, 17, 20, 3, 22, 26, 10, -4, 10, 11, 19, 17, 5, 15, 11, 10, 6, 7, 9, 8, -28, 8, 15, 21, 20, 9, 13, -5, 2, 0, -3, 8, 32, 27, -41, 4, 28, 12, 13, 4, 5, -16, -13, 7, -7, -18, 8, 24, -25, 13, 2, -6, -20, 0, -7, -11, -8, 22, 9, -9, 7, 30, -2, -20, -50, -37, -10, -6, 3, -12, -41, -8, -2, -11, 18, 9, -10, 6, -20, -34, -11, 0, 13, -17, -11, 5, 15, 20, 18, 2, -5, 4, 30, 8, -7, 3, -14, -20, 4, 4, 18, 29, 0, 2, 6, 7, 10, 17, 3, -2, 9, 9, 15, 0, 7, 23, -1, -1, -10, 32, -10, 16, 9, 19, 27, 37, 27, 1, 10, 21, 17, -5, 6, 5, -8, 16, 30, 32, 44, 41, 34, 24, -4, 13, 2, -16, -6, -10, -5, -14, -42, 13, -6, -31, -2, -12, -14, -4, 2, 9 },
{ -8, 5, 9, 29, 43, 32, 23, -22, 43, 56, 29, 21, -3, 4, 3, -21, 7, 24, 36, 42, 12, 7, 2, -2, 9, 9, 3, 3, 6, -17, 12, 8, 16, 5, 8, -4, 11, 6, 0, 12, -4, -13, 9, 27, 15, 8, 6, 3, -1, 3, -4, -9, -3, 1, 2, -18, 18, 24, 9, -21, -4, 11, -4, -6, -19, -8, 4, 14, -14, -32, 16, 0, 4, -16, -9, 10, -4, -24, -7, -3, 13, 12, -46, -63, 16, -8, -15, 1, 6, 17, -14, -22, 6, 6, 10, 50, 49, -23, 5, -14, 4, 17, 18, 13, 9, 18, 8, 21, 20, 46, 26, 44, 2, -12, -6, 14, 27, 20, 17, 18, 11, 14, 33, 17, 33, 21, 7, 4, 2, -6, 5, 13, 14, 2, 3, -6, 6, 7, 0, 14, 11, 12, 1, -9, 5, 19, 8, 7, -6, -21, -22, -17, -38, 0, -4, -2, -9, 5, -3, 6, 9, 15, -10, -27, -31, -25, -16, -11, 1, -5, 4, 8, 0, 5, 0, 14, -6, -55, -50, -32, -15, 3, 3, -22, -21, -10, -2, -12, -26, -22, -27, -45, -27, -4, -9, 1 },
{ -6, 2, -2, 20, -9, -9, -17, -1, 14, 8, 4, 16, -5, 8, 8, -4, 13, 11, -8, -22, -39, -54, -50, -30, -21, -16, -9, 2, 5, 15, 33, -3, -9, -30, -29, -30, -18, -5, -10, -6, -33, -9, 11, 25, 6, 12, 16, 4, 7, 6, 1, -5, -6, -15, -53, -22, 16, 20, 27, 30, 40, 37, 51, 23, -20, -16, 8, 15, -48, -8, 18, 21, 45, 42, 41, 41, 26, 7, 5, 7, -4, -2, -33, 9, 18, -12, -10, -17, -30, -46, -63, -16, 14, 8, -19, -20, 2, 41, 11, -19, -50, -47, -53, -14, -12, -1, 5, 11, 11, -3, 3, 28, -1, -20, -52, -25, -8, -10, -1, -1, -3, 9, 0, -1, 15, 32, 26, -10, -6, -7, -7, -1, -5, 9, 1, -4, -1, -7, -4, 42, 9, 5, 1, -2, -1, 0, 1, 6, -6, -8, -13, -6, 24, 27, -3, -23, -3, 25, 9, -2, -2, 7, 11, -6, -9, 2, 19, -15, -8, -9, 33, 21, -3, -19, -12, -14, 9, -1, 2, -13, 20, 6, 7, -15, -8, 13, 43, 19, 23, 35, 15, 41, 24, 22, -1, -1 },
{ 2, -3, 0, -6, 29, 0, 14, 5, -4, 18, -11, -14, -3, -7, 5, -3, 8, 16, -21, -8, 11, 24, 31, 18, 29, -8, 4, 5, 2, 11, 13, 13, 14, 6, 2, 23, 12, 21, 6, 3, 24, -15, 31, 15, 12, 14, 11, -19, -22, -12, -6, -4, -1, 5, 22, 47, 39, 5, 15, 16, -5, -22, 18, -5, -24, -2, 6, 14, 31, 7, 46, 22, -1, -6, -4, 15, 44, 9, 2, 4, 9, 6, 15, 8, 40, 14, 3, 11, 28, 33, 5, 6, 23, 5, -14, -16, -22, 2, 16, 0, 12, 16, 17, -15, -33, 6, 9, 9, 9, 22, -2, -30, 16, 12, 12, 18, -4, -31, -32, -7, -5, 8, 16, 20, -9, -42, 21, 29, 17, 8, 16, -18, -16, 10, 9, 10, 18, -1, -21, -27, 5, -9, -3, 7, 3, 7, -6, 19, 19, 14, 2, -16, -35, -23, -2, -18, -25, -21, -29, -14, -3, 30, 31, 23, -14, -45, -51, 19, 0, -3, 13, 5, -1, -3, 0, 20, 4, -15, -24, -44, -27, 21, 0, -13, -23, -6, 9, 6, 7, -8, 17, 1, -1, 24, -19, 0 },
{ -9, 3, 1, 34, 34, 49, 62, -22, -8, 37, 25, 22, -5, 2, 0, 4, 10, 2, 0, 25, 9, -5, -9, 26, 33, 65, 9, 9, -2, -36, -33, -10, 0, -1, 11, 2, 11, 16, 14, 17, 36, 29, -39, -31, -20, -12, -5, 2, 18, 25, 28, 10, 3, -1, 32, 1, -36, 2, -13, 1, 6, 5, 1, 4, -4, 3, -2, -22, 26, -4, -41, -37, 2, 18, 19, 10, 9, -20, -11, -6, -5, 7, 15, -18, -31, -16, -7, 17, 10, 10, 19, 3, 9, 11, 24, 38, 4, -53, -11, -45, -20, 0, 8, 28, 6, 5, 16, 31, 3, 6, -14, -43, -23, -35, -32, 10, 25, 32, -2, -14, 28, 7, 2, -7, -13, -42, -17, -37, 2, 5, 0, 19, -9, -2, 12, 0, -5, -14, -38, -29, 14, -39, -3, 8, 1, -4, 18, 19, -9, -12, -21, -3, -44, -23, -17, 1, -19, -7, 0, 20, 27, 22, 9, 2, -9, 0, -17, -20, 8, 0, -7, -12, -13, 7, 10, 16, 11, 13, -2, -10, -21, -26, -5, 4, 26, 5, -14, -4, -2, -9, 0, -15, -7, -26, 4, 8 },
{ -2, 7, -10, -25, -29, -23, -35, -34, -45, -25, -17, -7, 9, -4, -4, -25, -14, -44, -52, -23, -36, -27, -2, -20, 1, -19, -29, 0, -13, -14, -21, -13, -3, 9, -2, 3, 0, -5, 4, -6, -7, -23, -14, 16, 11, 8, 9, 5, -3, -21, -12, 10, -8, 13, -9, 10, 23, 14, 16, 3, 8, 8, 2, -33, 15, 16, -8, 4, 11, -12, 46, 5, 0, 1, 13, 18, 7, -61, 14, 24, 1, -12, -24, -16, 31, 6, -5, 10, 7, 29, 19, -67, 1, 23, 14, -4, -17, 10, -9, -3, 7, 22, 16, 24, -18, -41, 12, 19, 0, -5, -14, 3, -22, -13, 19, 11, 4, -9, -54, -6, 24, 11, 2, -15, -23, -21, 13, -5, 22, 1, -18, -46, -27, 16, 15, 6, -11, -14, -16, 13, -5, 11, -9, -20, -27, -9, 13, -1, 4, 1, -9, -7, -1, 21, -2, -5, -11, -10, -4, 11, 11, 5, 4, 3, 9, 9, 24, 5, 9, -10, -27, -8, -4, -2, 7, 3, 12, -4, 1, -8, -17, 3, 2, -5, -29, -23, -22, -18, -12, -22, -13, -10, -29, -6, -18, -1 },
{ 1, -7, -9, 5, -17, 1, -20, 12, 19, -2, 4, 4, 7, 8, -4, 21, 17, 33, 23, 10, 11, 5, 12, 19, 22, -17, 0, 2, 1, 27, 41, 16, 5, 0, 8, 7, 7, 3, 1, 9, 6, -12, 26, 34, 11, 2, 17, 22, 9, -2, 6, 8, 1, 1, -11, 11, 11, 3, 4, 7, 4, 10, 8, 1, 3, 0, -5, 10, -26, 5, -1, -4, -10, -3, -22, -32, -52, 1, -12, -20, -27, -18, -25, 7, 12, -17, -67, -83, -68, -60, -21, 16, 2, -3, -15, -28, 14, 44, -1, -23, -38, -23, -23, 2, 23, 30, 14, 19, 24, 20, 39, 32, 13, 22, 13, 26, 15, -1, 28, 5, 7, 19, 24, 20, 39, 49, -7, 40, 35, 31, 29, 10, 2, 10, 4, 4, 2, -6, 34, 45, -15, 44, 7, 17, 17, 0, 7, 16, 7, -2, -9, -3, 21, 14, 14, 10, 27, -5, -15, -4, -14, -10, 0, -7, -14, -9, -5, 35, 9, 33, 18, 7, 10, -1, 2, -1, -7, -29, -12, -21, 0, 13, 9, -4, -19, 9, 18, 21, -2, 17, 5, 9, 1, -29, 0, 1 },
{ 7, 0, 3, 18, 31, 49, 56, 47, 73, 34, 7, 17, -9, -7, 5, 18, 10, -6, -3, 4, 20, 23, 14, 39, 44, 24, 34, -2, -5, -13, -39, -16, -12, 16, 10, 14, 18, 25, 22, 38, 42, 39, 0, -17, -28, -1, 15, 21, 28, 31, 16, 14, 8, -9, 25, 31, 7, -19, -21, -7, 15, 32, 9, -24, -39, -57, -63, -77, -49, 18, -26, -15, -1, 17, 11, 3, -29, -24, 13, -15, -31, -49, -71, 3, -21, 2, 7, 13, -1, -12, -25, -7, 14, 28, 28, 32, -20, -23, -2, -21, -3, -2, -2, -2, -24, -17, 4, 8, 20, 20, 12, -39, -17, -4, -5, -15, -12, 0, -17, -18, 9, 17, 6, -2, 3, -47, -20, 9, 3, -4, -12, 0, -35, -2, 13, 0, 4, -2, 25, -38, -24, 3, 13, -2, 4, 5, 0, 16, 14, 2, 2, 5, 32, -17, -4, -7, 3, -7, 4, 5, 7, 14, 8, -3, 0, 6, 18, 16, -8, 4, 5, 2, -7, -9, 1, -6, 1, 4, 28, 25, 11, -12, 6, -5, -2, -10, 20, -14, 4, 19, 24, 32, 34, 20, 18, 4 },
{ -5, 4, 4, 19, 38, 42, 39, 23, 24, 46, 34, 19, 7, -8, -1, 13, 13, 35, 41, 37, 43, 33, 11, 12, 18, 35, -12, -7, -3, 2, 0, -5, -9, -9, -8, -10, -17, -17, -36, -35, -49, -34, -7, -30, -30, -14, -17, -7, 4, 18, 5, -13, -24, -47, -63, -67, 7, -10, -15, 0, 7, 4, 13, 42, -3, -20, -17, -27, -56, -35, 1, 14, 3, 17, 9, 10, 19, 11, -23, 9, 17, 9, -10, -39, -11, 24, 8, 11, 7, 4, 0, -8, -3, 4, 5, 21, 6, -42, -11, -16, 8, 9, 15, 16, 3, -6, -12, -6, 13, 9, 15, -41, 5, -26, 3, -5, 3, 31, -1, -12, -10, 10, 2, -4, 4, -10, 24, -21, -35, -28, -6, 6, 2, 11, -5, 11, 11, -1, 3, -3, 9, -18, -16, -21, -15, -3, 30, 21, -3, -4, -6, -17, 12, 14, 5, -12, -24, -34, -19, -9, 1, -7, -11, -27, -17, -1, -9, 5, -7, -7, 5, -16, 6, -6, -2, -16, -1, -2, 6, 6, 14, 14, 0, 12, 10, 15, 33, 35, 15, 33, 32, 17, 35, 11, 13, 0 },
{ -1, 9, -8, -9, -13, -19, -8, -8, 19, -46, -34, -17, 0, -9, 1, -6, -12, -38, -33, -21, -2, 5, 4, -15, -23, -11, 3, -2, -1, 0, -9, -1, -10, 4, 20, 28, 24, 15, 2, -20, 3, 3, 30, 25, 0, -5, 0, 16, 21, 24, 23, 17, 8, -1, -5, 1, 22, 18, -9, 5, 5, -2, -11, 2, 11, 32, 17, 15, -3, 9, 15, 32, 1, 2, -7, -34, -21, -6, -3, 28, 25, 9, -25, -7, 13, 17, 3, -11, -18, -16, -5, -13, -3, 25, 29, -7, -2, 17, 20, 0, -5, -2, -10, -1, 1, 9, 8, 17, 7, -5, -5, 24, 19, 9, -6, -8, 6, 2, -1, 0, 16, -6, -21, 6, -3, 21, 25, 12, 4, -5, 5, 2, -19, -2, 1, -8, -12, -12, -14, -13, 18, 8, 19, 22, 3, -14, -8, -5, -9, -15, -18, -20, -15, -4, -1, 4, -13, 22, 10, 5, 8, -1, -5, -7, -19, 2, 12, -20, 4, 14, 16, 30, 7, 21, 14, 18, 17, 5, -6, -20, 9, 6, 9, -9, -13, 27, 54, 31, 16, 17, 23, 39, 18, 2, -1, -1 },
{ -7, -8, -11, -14, -25, -30, -46, -13, -11, -30, -17, -7, -5, 0, -2, 4, -5, -4, 5, 3, 0, -27, -27, -63, -59, -43, -26, -9, 3, 38, 9, 9, 4, 23, 22, 6, -13, -26, -43, -35, -21, -17, 21, 43, 13, -1, -1, 8, 30, 25, 19, -12, -34, -61, -61, -5, 9, 16, 7, -11, 0, 1, -4, 41, 40, 13, -44, -75, -99, -5, 10, 39, 6, -10, -16, -13, -10, 28, 55, 26, -29, -69, -49, 11, 2, 27, -15, -16, -10, -7, 1, 28, 27, 9, -34, -46, 15, 43, 9, 28, -13, -10, 0, -11, -5, 15, 20, -8, -25, -6, 0, 41, 13, 13, -16, 0, 1, -14, 12, 17, 15, -10, 1, 20, 17, 57, 22, 16, -5, -10, -15, -4, -5, -8, -3, 1, 11, 7, 2, 35, 16, 22, -12, -14, -9, -8, -18, -18, -7, 3, 6, 1, 18, 16, 13, 27, 10, -4, -10, 3, -9, -10, -13, -3, 5, 6, 19, -11, -9, 2, 32, 13, -15, -10, -9, 6, 0, -7, 22, -2, 11, 26, 9, 9, 14, 22, 67, 38, 25, 29, 31, 33, 16, 11, 7, -7 },
{ -7, 0, -6, -2, 18, 7, -4, 15, -17, 26, -1, -12, 4, 8, -4, -7, -10, -7, -10, -9, -4, 16, 0, -8, -12, 2, -8, 7, 3, -2, -1, -15, -29, -18, -9, 8, 8, 12, 11, 9, 1, -4, -16, -19, -20, -44, -37, -17, -16, -2, -5, -3, 1, 6, 21, 22, -32, -28, -32, -26, -29, 0, 7, -7, -6, -11, -7, -16, -11, -9, -21, -49, -27, -13, 0, 6, -10, -5, -3, -23, -19, -50, -45, -8, -15, -20, -7, 9, 15, 16, 10, -1, 0, -7, -8, -17, -33, -17, -17, 16, 23, 15, 8, 0, 16, 30, 2, -25, -19, -25, -8, 36, -22, 21, 20, 11, 16, 5, 11, 26, -6, -19, -3, -9, 8, 41, -24, 17, 2, 4, 8, -13, 11, 16, 2, 5, 12, 7, 45, 25, -8, 19, 9, 9, 4, -8, -21, 6, 32, 36, 35, 24, 29, 9, -5, 6, 17, -2, -3, -10, -17, -4, 15, 33, 43, 8, -7, 11, -4, -32, -22, -15, -21, -11, -28, -23, -27, -17, 3, 10, -4, 25, -3, -13, -18, -38, -35, -25, -40, -40, -25, -33, -28, -30, -7, -7 },
{ 9, 3, -7, -12, -12, -11, 1, 17, -4, -30, -31, -18, -4, -1, -5, -16, -8, 8, -5, -2, 10, 21, 11, -19, -17, 4, 6, -4, 0, -6, 2, 2, -7, 2, 19, 17, 18, 22, 18, 6, 4, -3, -9, -23, 6, -2, 2, -6, -2, -3, -10, -3, -9, 0, -9, -11, -26, -3, -5, -8, -1, 6, 6, -11, -15, -8, 1, -8, -33, -11, -28, -6, 1, 2, -2, -4, -2, -15, 6, 1, -17, -27, -32, -31, -13, -16, -11, -7, -2, 3, 3, 2, 10, 5, 18, 11, 25, 5, -8, 7, -7, 2, 10, 16, 18, 20, 16, -4, -1, -6, 5, 62, -9, 17, -2, 2, 27, 19, 27, 34, 4, -7, 2, -4, 17, 38, -20, 13, 9, 6, 11, -12, -4, 17, 9, -1, 7, 20, 30, 34, -2, 29, 19, 23, 6, -7, -10, 16, 13, 13, 23, 29, 7, 15, 2, 11, 23, 13, 12, 0, -9, 13, 12, 18, 24, 24, -4, 1, -3, -45, -60, -44, -23, -10, -16, 3, 0, 9, 5, 0, -2, 12, 7, -17, 2, -23, -47, -38, -61, -72, -66, -69, -74, -36, -3, 1 },
{ 0, 5, -12, -14, 8, 7, 15, 27, 13, -33, -37, -7, -8, 9, -5, 11, -4, 13, 26, 50, 44, 36, 24, 17, -16, -9, 0, -7, 1, 12, -26, -5, -43, -67, -52, -28, -10, 15, 2, -14, -21, 0, -5, 2, -23, -39, -96, -86, -29, 17, 29, 36, 25, -9, -30, -12, -23, -6, -41, -68, -39, -4, -1, -8, 5, 9, 6, 23, -16, -6, -13, -16, -37, -22, 5, -1, -36, -31, 2, 10, 11, 3, -7, 6, -30, -10, -23, -5, 3, -1, -24, 23, 17, 26, 17, 6, 13, 19, -16, -25, 1, -2, -4, 5, 14, 22, 20, 2, -8, -28, -11, 24, 23, -13, 4, 14, 10, 21, 22, -1, 0, -12, -28, -24, 1, 10, 8, -1, -4, -5, 10, 2, -1, 2, -2, 3, 6, 16, 18, 21, 2, 9, 26, 2, -13, -19, 3, 2, -2, -1, -16, 11, 19, -22, 3, 13, 6, -1, -10, -24, -21, -10, -14, -16, -17, -10, -23, -12, -7, -11, 10, 4, 6, -12, 0, 6, 3, 0, 5, 3, -27, -3, 6, 14, 14, 34, 25, 28, 29, 58, 56, 50, 70, 6, -22, 2 },
{ -5, -6, 6, 27, 32, 46, 29, -14, 3, 40, 39, 29, 2, 9, -6, 5, 16, 31, 16, 21, 23, 21, 3, 17, 25, 6, -3, -4, -1, 9, 20, 20, 13, 0, -13, -15, -21, -15, -15, -28, -19, -39, 6, 13, 10, 7, 20, 1, 7, 10, 9, -18, -15, -5, -13, 10, -14, 24, 5, 3, -1, -20, -1, 3, -6, -15, -11, -9, -30, -15, -5, 12, -19, -4, -15, -10, 5, -5, 4, 9, 4, -24, -61, -38, 3, -3, -29, 8, 2, 20, 11, 11, 25, 28, 25, 5, -38, -37, -4, 7, -11, -8, 5, 23, 14, 1, 28, 21, 23, -8, -61, -41, 25, -19, -50, -32, 2, 25, 0, 12, 15, 1, 1, -2, -41, -29, -15, 25, -8, -28, -43, -1, 10, 7, 6, -8, -19, -28, -51, 15, 6, 37, -16, -11, -20, -18, 3, 2, 3, -18, -30, -41, -17, -10, -5, 15, -9, -4, 9, 5, -7, -10, -11, -12, -27, -18, -17, 18, 1, 29, 33, 28, 20, 11, -4, -13, -6, -3, 0, -17, -22, 1, -1, 15, 44, 46, 38, 23, 9, 10, 18, 14, 0, -3, 6, 5 }
};


wire dense1_en = enable;
    reg dense1_terminat;

    
    dense_layer #(.numar_neuroni(32),.dimensiune_intrare(196), .latime(8)) dense_layer1(.clock(clock), .layer_enable(dense1_en), .reset(reset),
                                                                        .date_intrare(imagine_trasa), .weights(VECTOR_WEIGHTS_LAYER2), .biases(VECTOR_BIASURI_LAYER2),
                                                                        .date_iesire(dense1_retea), .layer_terminat(dense1_terminat)); //Dense layer
    
    relu relu_activation[31:0] (.date_intrare(dense1_retea), .date_iesire(relu_retea)); 
    assign iesire_layer = relu_retea;               
    assign layer_terminat = dense1_terminat;

endmodule